library verilog;
use verilog.vl_types.all;
entity pipelinedProc_vlg_vec_tst is
end pipelinedProc_vlg_vec_tst;
